
module Decoder(
	n_T0, n_T1X,
	n_T2, n_T3, n_T4, n_T5, 
	IR01,
	IR, n_IR,
	X);

	input n_T0;
	input n_T1X;
	input n_T2;
	input n_T3;
	input n_T4;
	input n_T5; 
	input IR01;
	input [7:0] IR;
	input [7:0] n_IR;

	output [129:0] X;

	wire [20:0] d;
	assign d = {n_T1X,n_T0,n_IR[5],IR[5],n_IR[6],IR[6],n_IR[2],IR[2],n_IR[3],IR[3],n_IR[4],IR[4],n_IR[7],IR[7],n_IR[0],IR01,n_IR[1],n_T2,n_T3,n_T4,n_T5};

	assign X[0] = ~|{d[5],d[8],d[14],d[15],d[17]};
	assign X[1] = ~|{d[2],d[6],d[10],d[11],d[13]};
	assign X[2] = ~|{d[3],d[6],d[10],d[12],d[13]};
	assign X[3] = ~|{d[5],d[8],d[9],d[12],d[13],d[17],d[19]};
	assign X[4] = ~|{d[5],d[8],d[10],d[12],d[13],d[15],d[17],d[19]};
	assign X[5] = ~|{d[5],d[8],d[9],d[16],d[17],d[19]};
	assign X[6] = ~|{d[3],d[10],d[14]};
	assign X[7] = ~|{d[4],d[8],d[15]};
	assign X[8] = ~|{d[3],d[6],d[9],d[11],d[13]};
	assign X[9] = ~|{d[4],d[8],d[9],d[12],d[13],d[15],d[17],d[19]};
	assign X[10] = ~|{d[4],d[8],d[9],d[12],d[13],d[16],d[17],d[19]};
	assign X[11] = ~|{d[5],d[8],d[9],d[16],d[18],d[19]};
	assign X[12] = ~|{d[4],d[8],d[15],d[17]};
	assign X[13] = ~|{d[4],d[8],d[10],d[12],d[13],d[15],d[17],d[19]};
	assign X[14] = ~|{d[4],d[8],d[15],d[18],d[19]};
	assign X[15] = ~|{d[4],d[8],d[9],d[12],d[13],d[16],d[17],d[20]};
	assign X[16] = ~|{d[5],d[8],d[9],d[12],d[13],d[16],d[18],d[20]};
	assign X[17] = ~|{d[4],d[8],d[10],d[12],d[13],d[15],d[18],d[19]};
	assign X[18] = ~|{d[5],d[8],d[9],d[12],d[13],d[17],d[20]};
	assign X[19] = ~|{d[5],d[8],d[14],d[15],d[18],d[19]};
	assign X[20] = ~|{d[5],d[8],d[9],d[15],d[18],d[19]};
	assign X[21] = ~|{d[5],d[7],d[9],d[11],d[13],d[15],d[18],d[19]};
	assign X[22] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[15],d[17]};
	assign X[23] = ~|{d[5],d[7],d[9],d[12],d[13],d[17],d[19]};
	assign X[24] = ~|{d[1],d[5],d[7],d[9],d[11],d[13],d[16],d[18]};
	assign X[25] = ~|{d[2],d[5],d[7],d[9],d[12],d[13],d[18]};
	assign X[26] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[16],d[17]};
	assign X[27] = ~|{d[4],d[7],d[16],d[18]};
	assign X[28] = ~|{d[3]};
	assign X[29] = ~|{d[6],d[7],d[16],d[17],d[19]};
	assign X[30] = ~|{d[5],d[7],d[9],d[12],d[14],d[16]};
	assign X[31] = ~|{d[3],d[9],d[12],d[14]};
	assign X[32] = ~|{d[6],d[7],d[15],d[17],d[19]};
	assign X[33] = ~|{d[3],d[11]};
	assign X[34] = ~|{d[19]};
	assign X[35] = ~|{d[3],d[5],d[7],d[9],d[13]};
	assign X[36] = ~|{d[2],d[5],d[7],d[9]};
	assign X[37] = ~|{d[1],d[5],d[7],d[9],d[11],d[13],d[15]};
	assign X[38] = ~|{d[1],d[5],d[7],d[9],d[11],d[13],d[16],d[17]};
	assign X[39] = ~|{d[2],d[6],d[9],d[11],d[13]};
	assign X[40] = ~|{d[1],d[6],d[10],d[11],d[13]};
	assign X[41] = ~|{d[3],d[6],d[10],d[11],d[13]};
	assign X[42] = ~|{d[2],d[10],d[12]};
	assign X[43] = ~|{d[5],d[7],d[9],d[12],d[13],d[18]};
	assign X[44] = ~|{d[4],d[8],d[16],d[18]};
	assign X[45] = ~|{d[1],d[6],d[9],d[11],d[13]};
	assign X[46] = ~|{d[2],d[6],d[10],d[11],d[13]};
	assign X[47] = ~|{d[5],d[7],d[9],d[11],d[13],d[16]};
	assign X[48] = ~|{d[3],d[5],d[7],d[9],d[11],d[13],d[15],d[18]};
	assign X[49] = ~|{d[5],d[8],d[9],d[16],d[19]};
	assign X[50] = ~|{d[6],d[8],d[16],d[17],d[19]};
	assign X[51] = ~|{d[6],d[8],d[16],d[18],d[19]};
	assign X[52] = ~|{d[6],d[16],d[18],d[19]};
	assign X[53] = ~|{d[4],d[7],d[15],d[18]};
	assign X[54] = ~|{d[2],d[5],d[7],d[9],d[12],d[14],d[16]};
	assign X[55] = ~|{d[4],d[7],d[15]};
	assign X[56] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[15],d[18]};
	assign X[57] = ~|{d[3],d[5],d[7],d[9],d[13]};
	assign X[58] = ~|{d[5],d[8],d[10],d[12],d[13],d[15],d[17],d[19]};
	assign X[59] = ~|{d[6],d[7],d[20]};
	assign X[60] = ~|{d[6],d[16],d[18],d[20]};
	assign X[61] = ~|{d[4],d[7],d[9],d[12],d[13],d[20]};
	assign X[62] = ~|{d[4],d[8],d[9],d[12],d[13],d[15],d[17],d[19]};
	assign X[63] = ~|{d[5],d[7],d[9],d[12],d[13],d[16],d[18],d[19]};
	assign X[64] = ~|{d[6],d[8],d[15],d[18],d[19]};
	assign X[65] = ~|{d[6],d[19]};
	assign X[66] = ~|{d[5],d[8],d[9],d[12],d[13],d[15],d[18],d[19]};
	assign X[67] = ~|{d[4],d[7],d[9],d[12],d[13],d[19]};
	assign X[68] = ~|{d[4],d[8],d[9],d[12],d[13],d[15],d[18],d[19]};
	assign X[69] = ~|{d[5],d[7],d[9],d[14],d[15],d[18],d[19]};
	assign X[70] = ~|{d[6],d[7],d[15],d[18],d[19]};
	assign X[71] = ~|{d[1],d[10],d[12]};
	assign X[72] = ~|{d[0],d[6],d[10],d[11],d[13]};
	assign X[73] = ~|{d[5],d[10],d[11],d[13],d[19]};
	assign X[74] = ~|{d[3],d[5],d[7],d[9],d[12],d[13],d[16],d[17]};
	assign X[75] = ~|{d[4],d[7],d[9],d[12],d[13],d[16],d[19]};
	assign X[76] = ~|{d[4],d[7],d[16]};
	assign X[77] = ~|{d[3],d[5],d[7],d[9],d[11],d[13],d[15],d[17]};
	assign X[78] = ~|{d[2],d[5],d[7],d[9],d[11],d[13],d[15],d[18]};
	assign X[79] = ~|{d[6],d[8],d[15],d[17]};
	assign X[80] = ~|{d[3],d[5],d[10],d[11],d[13]};
	assign X[81] = ~|{d[3],d[11],d[14]};
	assign X[82] = ~|{d[3],d[6],d[11],d[13]};
	assign X[83] = ~|{d[3],d[12]};
	assign X[84] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[16],d[18]};
	assign X[85] = ~|{d[1]};
	assign X[86] = ~|{d[2]};
	assign X[87] = ~|{d[5],d[7],d[9],d[11],d[13],d[17],d[19]};
	assign X[88] = ~|{d[5],d[7],d[9],d[12],d[14],d[16],d[19]};
	assign X[89] = ~|{d[0],d[6],d[9],d[11],d[13]};
	assign X[90] = ~|{d[2],d[12]};
	assign X[91] = ~|{d[1],d[6],d[10],d[11],d[13]};
	assign X[92] = ~|{d[2],d[10],d[12]};
	assign X[93] = ~|{d[2],d[5],d[10],d[11],d[13]};
	assign X[94] = ~|{d[5],d[7],d[9],d[11],d[13],d[17]};
	assign X[95] = ~|{d[5],d[7],d[9],d[11],d[13],d[15],d[18]};
	assign X[96] = ~|{d[5],d[7],d[9],d[12],d[14],d[16]};
	assign X[97] = ~|{d[8],d[15],d[17]};
	assign X[98] = ~|{d[1],d[5],d[7],d[9],d[11],d[13],d[15],d[17]};
	assign X[99] = ~|{d[3],d[5],d[7],d[9],d[12],d[13],d[15],d[17]};
	assign X[100] = ~|{d[3],d[5],d[7],d[9],d[12],d[13],d[17]};
	assign X[101] = ~|{d[1],d[5],d[7],d[9],d[12],d[14],d[16]};
	assign X[102] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[16]};
	assign X[103] = ~|{d[0],d[5],d[7],d[9],d[11],d[13],d[15],d[18]};
	assign X[104] = ~|{d[3],d[5],d[7],d[9],d[12],d[14],d[16],d[17]};
	assign X[105] = ~|{d[2],d[5],d[7],d[9],d[12],d[13],d[18]};
	assign X[106] = ~|{d[4],d[16]};
	assign X[107] = ~|{d[4],d[7],d[15]};
	assign X[108] = ~|{d[5],d[7],d[10],d[12],d[13],d[16],d[19]};
	assign X[109] = ~|{d[5],d[7],d[9],d[14],d[15],d[18],d[20]};
	assign X[110] = ~|{d[5],d[7],d[10],d[12],d[13],d[15],d[19]};
	assign X[111] = ~|{d[2],d[10],d[11],d[14]};
	assign X[112] = ~|{d[6],d[16],d[18],d[20]};
	assign X[113] = ~|{d[5],d[7],d[9],d[14],d[15],d[18],d[19]};
	assign X[114] = ~|{d[5],d[7],d[9],d[12],d[13],d[15],d[18],d[19]};
	assign X[115] = ~|{d[1],d[5],d[7],d[9],d[11],d[13],d[16],d[17]};
	assign X[116] = ~|{d[6],d[8],d[16],d[17],d[20]};
	assign X[117] = ~|{d[5],d[8],d[9],d[12],d[14],d[16],d[20]};
	assign X[118] = ~|{d[4],d[7],d[9],d[12],d[13],d[15],d[20]};
	assign X[119] = ~|{d[5],d[8],d[9],d[11],d[16],d[20]};
	assign X[120] = ~|{d[5],d[8],d[10],d[12],d[13],d[16],d[19]};
	assign X[121] = ~|{d[15]};
	assign X[122] = ~|{d[2],d[9],d[12],d[14]};
	assign X[123] = ~|{d[3],d[9],d[11],d[14]};
	assign X[124] = ~|{d[0],d[6],d[11],d[13]};
	assign X[125] = ~|{d[1],d[10],d[12]};
	assign X[126] = ~|{d[7]};
	assign X[127] = ~|{d[5],d[8],d[10],d[12],d[13],d[15],d[18]};
	assign X[128] = ~|{d[12],d[13]};
	assign X[129] = ~|{d[5],d[7],d[9],d[12],d[13]};

endmodule // Decoder
