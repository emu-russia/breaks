
module PixelClock(
	n_CLK, CLK, RES,
	n_PCLK, PCLK);

	input n_CLK;
	input CLK;
	input RES;

	output n_PCLK;
	output PCLK;

endmodule // PixelClock
