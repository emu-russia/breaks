// Тестовая программа на Verilog

// Пока мы модули не используем, будем считать что мы уже внутри модуля.
//module test;

    // балуемся с числами (пока просто поток токенов, парсера всё равно нет)
    123     // десятичное
    0234    // с нуля
    01_22_33    // с черточками

    8 'b 11001100   // двоичное 8 разрядов
    8 'b ?1x0_Z1z0   // двоичное 8 разрядов, с черточками и пр.
    4 'b 10012      // ошибка! цифра 2

    2 'o 35
    2 'o 35_22
    2 'o 35_28      // ошибка! цифра 8

    2 'h 1234_5678_ab
    2 'h 35_G       // G!
    2 'h 00035_28 
    

    parameter DUMMY = 1, NBIT = 4;
    input CLK;

    wire a, b, c;
    wire [7:0] ___busa;
    wire [0:9] busb;
    wand vectored [7:0] andbus;
    reg [NBIT-1:0] dout;
    trireg [7:0] treg;

    reg MYREG2;

    always @ (CLK)
        MYREG2 = MYREG2 ^ 1;
    end

//endmodule
