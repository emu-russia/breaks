
module ClkGen(PHI0, PHI1, PHI2, PHI1_topad, PHI2_topad);

	input PHI0;
	output PHI1;
	output PHI2;
	output PHI1_topad;
	output PHI2_topad;

endmodule 	// ClkGen
