
module ExtraCounter(
	PHI1, PHI2, TRES2, n_ready, T1,
	n_T2, n_T3, n_T4, n_T5);

	input PHI1;
	input PHI2;
	input TRES2;
	input n_ready;
	input T1;

	output n_T2;
	output n_T3;
	output n_T4;
	output n_T5;

endmodule // ExtraCounter
